module multiplier_19_bits
	#(
		parameter d_width = 20
	)
	(
		input [d_width-1:0] A ,
		input [d_width-1:0] B ,
		output [2*d_width-1:0] mul
	);
	
	// generate partial products
	wire [d_width-1:0] pp [d_width-1:0] ;
	
	genvar i;
   generate
   for (i = 0; i < 19; i=i+1) begin:n
		 assign pp[0][i] = A[i] & B[0] ;
		 assign pp[1][i] = A[i] & B[1] ;
		 assign pp[2][i] = A[i] & B[2] ;
		 assign pp[3][i] = A[i] & B[3] ;
		 assign pp[4][i] = A[i] & B[4] ;
		 assign pp[5][i] = A[i] & B[5] ;
		 assign pp[6][i] = A[i] & B[6] ;
		 assign pp[7][i] = A[i] & B[7] ;
		 assign pp[8][i] = A[i] & B[8] ;
		 assign pp[9][i] = A[i] & B[9] ;
		 assign pp[10][i] = A[i] & B[10] ;
		 assign pp[11][i] = A[i] & B[11] ;
		 assign pp[12][i] = A[i] & B[12] ;
		 assign pp[13][i] = A[i] & B[13] ;
		 assign pp[14][i] = A[i] & B[14] ;
		 assign pp[15][i] = A[i] & B[15] ;
		 assign pp[16][i] = A[i] & B[16] ;
		 assign pp[17][i] = A[i] & B[17] ;
		 assign pp[18][i] = A[i] & B[18] ;
	end
	endgenerate
	
	// level-7, capacity-19, lines -37, our max bit length size of line size-19
	wire       l7_line1 ;
   wire [1:0] l7_line2 ;
   wire [2:0] l7_line3 ;
   wire [3:0] l7_line4 ;
   wire [4:0] l7_line5 ;
   wire [5:0] l7_line6 ;
   wire [6:0] l7_line7 ;
   wire [7:0] l7_line8 ;
   wire [8:0] l7_line9 ;
   wire [9:0] l7_line10 ;
   wire [10:0] l7_line11 ;
   wire [11:0] l7_line12 ;
   wire [12:0] l7_line13 ;
   wire [13:0] l7_line14 ;
   wire [14:0] l7_line15 ;
   wire [15:0] l7_line16 ;
   wire [16:0] l7_line17 ;
   wire [17:0] l7_line18 ;
   wire [18:0] l7_line19 ;
	
	wire [17:0] l7_line20 ;
   wire [16:0] l7_line21 ;
   wire [15:0] l7_line22 ;
   wire [14:0] l7_line23 ;
   wire [13:0] l7_line24 ;
   wire [12:0] l7_line25 ;
   wire [11:0] l7_line26 ;
   wire [10:0] l7_line27 ;
   wire [9:0] l7_line28 ;
   wire [8:0] l7_line29 ;
   wire [7:0] l7_line30 ;
   wire [6:0] l7_line31 ;
   wire [5:0] l7_line32 ;
   wire [4:0] l7_line33 ;
   wire [3:0] l7_line34 ;
   wire [2:0] l7_line35 ;
   wire [1:0] l7_line36 ;
   wire       l7_line37 ;
	
	assign l7_line1 = { pp[0][0] };
   assign l7_line2 = { pp[1][0] , pp[0][1] };
   assign l7_line3 = { pp[2][0] , pp[1][1] , pp[0][2] };
   assign l7_line4 = { pp[3][0] , pp[2][1] , pp[1][2] , pp[0][3] };
   assign l7_line5 = { pp[4][0] , pp[3][1] , pp[2][2] , pp[1][3] , pp[0][4] };
   assign l7_line6 = { pp[5][0] , pp[4][1] , pp[3][2] , pp[2][3] , pp[1][4] , pp[0][5] };
   assign l7_line7 = { pp[6][0] , pp[5][1] , pp[4][2] , pp[3][3] , pp[2][4] , pp[1][5] , pp[0][6] };
   assign l7_line8 = { pp[7][0] , pp[6][1] , pp[5][2] , pp[4][3] , pp[3][4] , pp[2][5] , pp[1][6] , pp[0][7] };
   assign l7_line9 = { pp[8][0] , pp[7][1] , pp[6][2] , pp[5][3] , pp[4][4] , pp[3][5] , pp[2][6] , pp[1][7] , pp[0][8] };
   assign l7_line10 = { pp[9][0] , pp[8][1] , pp[7][2] , pp[6][3] , pp[5][4] , pp[4][5] , pp[3][6] , pp[2][7] , pp[1][8] , pp[0][9] };
   assign l7_line11 = { pp[10][0] , pp[9][1] , pp[8][2] , pp[7][3] , pp[6][4] , pp[5][5] , pp[4][6] , pp[3][7] , pp[2][8] , pp[1][9] , pp[0][10] };
   assign l7_line12 = { pp[11][0] , pp[10][1] , pp[9][2] , pp[8][3] , pp[7][4] , pp[6][5] , pp[5][6] , pp[4][7] , pp[3][8] , pp[2][9] , pp[1][10] , pp[0][11] };
   assign l7_line13 = { pp[12][0] , pp[11][1] , pp[10][2] , pp[9][3] , pp[8][4] , pp[7][5] , pp[6][6] , pp[5][7] , pp[4][8] , pp[3][9] , pp[2][10] , pp[1][11] , pp[0][12] };
   assign l7_line14 = { pp[13][0] , pp[12][1] , pp[11][2] , pp[10][3] , pp[9][4] , pp[8][5] , pp[7][6] , pp[6][7] , pp[5][8] , pp[4][9] , pp[3][10] , pp[2][11] , pp[1][12] , pp[0][13] };
   assign l7_line15 = { pp[14][0] , pp[13][1] , pp[12][2] , pp[11][3] , pp[10][4] , pp[9][5] , pp[8][6] , pp[7][7] , pp[6][8] , pp[5][9] , pp[4][10] , pp[3][11] , pp[2][12] , pp[1][13] , pp[0][14] };
   assign l7_line16 = { pp[15][0] , pp[14][1] , pp[13][2] , pp[12][3] , pp[11][4] , pp[10][5] , pp[9][6] , pp[8][7] , pp[7][8] , pp[6][9] , pp[5][10] , pp[4][11] , pp[3][12] , pp[2][13] , pp[1][14] , pp[0][15] };
   assign l7_line17 = { pp[16][0] , pp[15][1] , pp[14][2] , pp[13][3] , pp[12][4] , pp[11][5] , pp[10][6] , pp[9][7] , pp[8][8] , pp[7][9] , pp[6][10] , pp[5][11] , pp[4][12] , pp[3][13] , pp[2][14] , pp[1][15] , pp[0][16] };
   assign l7_line18 = { pp[17][0] , pp[16][1] , pp[15][2] , pp[14][3] , pp[13][4] , pp[12][5] , pp[11][6] , pp[10][7] , pp[9][8] , pp[8][9] , pp[7][10] , pp[6][11] , pp[5][12] , pp[4][13] , pp[3][14] , pp[2][15] , pp[1][16] , pp[0][17] };
   assign l7_line19 = { pp[18][0] , pp[17][1] , pp[16][2] , pp[15][3] , pp[14][4] , pp[13][5] , pp[12][6] , pp[11][7] , pp[10][8] , pp[9][9] , pp[8][10] , pp[7][11] , pp[6][12] , pp[5][13] , pp[4][14] , pp[3][15] , pp[2][16] , pp[1][17] , pp[0][18] };

	assign l7_line20 = { pp[18][1] , pp[17][2] , pp[16][3] , pp[15][4] , pp[14][5] , pp[13][6] , pp[12][7] , pp[11][8] , pp[10][9] , pp[9][10] , pp[8][11] , pp[7][12] , pp[6][13] , pp[5][14] , pp[4][15] , pp[3][16] , pp[2][17] , pp[1][18] };
   assign l7_line21 = { pp[18][2] , pp[17][3] , pp[16][4] , pp[15][5] , pp[14][6] , pp[13][7] , pp[12][8] , pp[11][9] , pp[10][10] , pp[9][11] , pp[8][12] , pp[7][13] , pp[6][14] , pp[5][15] , pp[4][16] , pp[3][17] , pp[2][18] };
   assign l7_line22 = { pp[18][3] , pp[17][4] , pp[16][5] , pp[15][6] , pp[14][7] , pp[13][8] , pp[12][9] , pp[11][10] , pp[10][11] , pp[9][12] , pp[8][13] , pp[7][14] , pp[6][15] , pp[5][16] , pp[4][17] , pp[3][18] };
   assign l7_line23 = { pp[18][4] , pp[17][5] , pp[16][6] , pp[15][7] , pp[14][8] , pp[13][9] , pp[12][10] , pp[11][11] , pp[10][12] , pp[9][13] , pp[8][14] , pp[7][15] , pp[6][16] , pp[5][17] , pp[4][18] };
   assign l7_line24 = { pp[18][5] , pp[17][6] , pp[16][7] , pp[15][8] , pp[14][9] , pp[13][10] , pp[12][11] , pp[11][12] , pp[10][13] , pp[9][14] , pp[8][15] , pp[7][16] , pp[6][17] , pp[5][18] };
   assign l7_line25 = { pp[18][6] , pp[17][7] , pp[16][8] , pp[15][9] , pp[14][10] , pp[13][11] , pp[12][12] , pp[11][13] , pp[10][14] , pp[9][15] , pp[8][16] , pp[7][17] , pp[6][18] };
   assign l7_line26 = { pp[18][7] , pp[17][8] , pp[16][9] , pp[15][10] , pp[14][11] , pp[13][12] , pp[12][13] , pp[11][14] , pp[10][15] , pp[9][16] , pp[8][17] , pp[7][18] };
   assign l7_line27 = { pp[18][8] , pp[17][9] , pp[16][10] , pp[15][11] , pp[14][12] , pp[13][13] , pp[12][14] , pp[11][15] , pp[10][16] , pp[9][17] , pp[8][18] };
   assign l7_line28 = { pp[18][9] , pp[17][10] , pp[16][11] , pp[15][12] , pp[14][13] , pp[13][14] , pp[12][15] , pp[11][16] , pp[10][17] , pp[9][18] };
   assign l7_line29 = { pp[18][10] , pp[17][11] , pp[16][12] , pp[15][13] , pp[14][14] , pp[13][15] , pp[12][16] , pp[11][17] , pp[10][18] };
   assign l7_line30 = { pp[18][11] , pp[17][12] , pp[16][13] , pp[15][14] , pp[14][15] , pp[13][16] , pp[12][17] , pp[11][18] };
   assign l7_line31 = { pp[18][12] , pp[17][13] , pp[16][14] , pp[15][15] , pp[14][16] , pp[13][17] , pp[12][18] };
   assign l7_line32 = { pp[18][13] , pp[17][14] , pp[16][15] , pp[15][16] , pp[14][17] , pp[13][18] };
   assign l7_line33 = { pp[18][14] , pp[17][15] , pp[16][16] , pp[15][17] , pp[14][18] };
   assign l7_line34 = { pp[18][15] , pp[17][16] , pp[16][17] , pp[15][18] };
   assign l7_line35 = { pp[18][16] , pp[17][17] , pp[16][18] };
   assign l7_line36 = { pp[18][17] , pp[17][18] };
   assign l7_line37 = { pp[18][18] };
	
	// partial product values put in lines... Now we have to reduce these lines...
	// for that Full Adders will be used
	// so, first next level lines have to be declared
	
	wire       l6_line1 ;
   wire [1:0] l6_line2 ;
   wire [2:0] l6_line3 ;
   wire [3:0] l6_line4 ;
   wire [4:0] l6_line5 ;
   wire [5:0] l6_line6 ;
   wire [6:0] l6_line7 ;
   wire [7:0] l6_line8 ;
   wire [8:0] l6_line9 ;
   wire [9:0] l6_line10 ;
   wire [10:0] l6_line11 ;
   wire [11:0] l6_line12 ;
   wire [12:0] l6_line13 ;
	
	wire [12:0] l6_line14 ;
   wire [12:0] l6_line15 ;
   wire [12:0] l6_line16 ;
   wire [12:0] l6_line17 ;
   wire [12:0] l6_line18 ;
   wire [12:0] l6_line19 ;
   wire [12:0] l6_line20 ;
   wire [12:0] l6_line21 ;
   wire [12:0] l6_line22 ;
   wire [12:0] l6_line23 ;
   wire [12:0] l6_line24 ;
   wire [12:0] l6_line25 ;
   wire [12:0] l6_line26 ;
	
	wire [10:0] l6_line27 ;
   wire [9:0] l6_line28 ;
   wire [8:0] l6_line29 ;
   wire [7:0] l6_line30 ;
   wire [6:0] l6_line31 ;
   wire [5:0] l6_line32 ;
   wire [4:0] l6_line33 ;
   wire [3:0] l6_line34 ;
   wire [2:0] l6_line35 ;
   wire [1:0] l6_line36 ;
   wire [0:0] l6_line37 ;
	
	// instantiating ful adders for level-6 in level-7
	HA level7_line14_HA1 ( l7_line14[0], l7_line14[1],              l6_line14[0], l6_line15[0]) ;
	
   FA level7_line15_FA1 ( l7_line15[0], l7_line15[1], l7_line15[2], l6_line15[1], l6_line16[0]) ;
   HA level7_line15_HA1 ( l7_line15[3], l7_line15[4],              l6_line15[2], l6_line16[1]) ;

   FA level7_line16_FA1 ( l7_line16[0], l7_line16[1], l7_line16[2], l6_line16[2], l6_line17[0]) ;
   FA level7_line16_FA2 ( l7_line16[3], l7_line16[4], l7_line16[5], l6_line16[3], l6_line17[1]) ;
   HA level7_line16_HA1 ( l7_line16[6], l7_line16[7],              l6_line16[4], l6_line17[2]) ;

   FA level7_line17_FA1 ( l7_line17[0], l7_line17[1], l7_line17[2], l6_line17[3], l6_line18[0]) ;
   FA level7_line17_FA2 ( l7_line17[3], l7_line17[4], l7_line17[5], l6_line17[4], l6_line18[1]) ;
   FA level7_line17_FA3 ( l7_line17[6], l7_line17[7], l7_line17[8], l6_line17[5], l6_line18[2]) ;
   HA level7_line17_HA1 ( l7_line17[9], l7_line17[10],              l6_line17[6], l6_line18[3]) ;

   FA level7_line18_FA1 ( l7_line18[0], l7_line18[1], l7_line18[2], l6_line18[4], l6_line19[0]) ;
   FA level7_line18_FA2 ( l7_line18[3], l7_line18[4], l7_line18[5], l6_line18[5], l6_line19[1]) ;
   FA level7_line18_FA3 ( l7_line18[6], l7_line18[7], l7_line18[8], l6_line18[6], l6_line19[2]) ;
   FA level7_line18_FA4 ( l7_line18[9], l7_line18[10], l7_line18[11], l6_line18[7], l6_line19[3]) ;
   HA level7_line18_HA1 ( l7_line18[12], l7_line18[13],              l6_line18[8], l6_line19[4]) ;

   FA level7_line19_FA1 ( l7_line19[0], l7_line19[1], l7_line19[2], l6_line19[5], l6_line20[0]) ;
   FA level7_line19_FA2 ( l7_line19[3], l7_line19[4], l7_line19[5], l6_line19[6], l6_line20[1]) ;
   FA level7_line19_FA3 ( l7_line19[6], l7_line19[7], l7_line19[8], l6_line19[7], l6_line20[2]) ;
   FA level7_line19_FA4 ( l7_line19[9], l7_line19[10], l7_line19[11], l6_line19[8], l6_line20[3]) ;
   FA level7_line19_FA5 ( l7_line19[12], l7_line19[13], l7_line19[14], l6_line19[9], l6_line20[4]) ;
   HA level7_line19_HA1 ( l7_line19[15], l7_line19[16],              l6_line19[10], l6_line20[5]) ;
	
	assign l6_line14[12:1] = l7_line14[13:2] ;
   assign l6_line15[12:3] = l7_line15[14:5] ;
   assign l6_line16[12:5] = l7_line16[15:8] ;
   assign l6_line17[12:7] = l7_line17[16:11] ;
   assign l6_line18[12:9] = l7_line18[17:14] ;
   assign l6_line19[12:11] = l7_line19[18:17] ;
	
	FA level7_line20_FA1 ( l7_line20[0], l7_line20[1], l7_line20[2], l6_line20[6], l6_line21[0]) ;
   FA level7_line20_FA2 ( l7_line20[3], l7_line20[4], l7_line20[5], l6_line20[7], l6_line21[1]) ;
   FA level7_line20_FA3 ( l7_line20[6], l7_line20[7], l7_line20[8], l6_line20[8], l6_line21[2]) ;
   FA level7_line20_FA4 ( l7_line20[9], l7_line20[10], l7_line20[11], l6_line20[9], l6_line21[3]) ;
   FA level7_line20_FA5 ( l7_line20[12], l7_line20[13], l7_line20[14], l6_line20[10], l6_line21[4]) ;
   HA level7_line20_HA1 ( l7_line20[15], l7_line20[16],              l6_line20[11], l6_line21[5]) ;
	
   FA level7_line21_FA1 ( l7_line21[0], l7_line21[1], l7_line21[2], l6_line21[6], l6_line22[0]) ;
   FA level7_line21_FA2 ( l7_line21[3], l7_line21[4], l7_line21[5], l6_line21[7], l6_line22[1]) ;
   FA level7_line21_FA3 ( l7_line21[6], l7_line21[7], l7_line21[8], l6_line21[8], l6_line22[2]) ;
   FA level7_line21_FA4 ( l7_line21[9], l7_line21[10], l7_line21[11], l6_line21[9], l6_line22[3]) ;
   FA level7_line21_FA5 ( l7_line21[12], l7_line21[13], l7_line21[14], l6_line21[10], l6_line22[4]) ;

   FA level7_line22_FA1 ( l7_line22[0], l7_line22[1], l7_line22[2], l6_line22[5], l6_line23[0]) ;
   FA level7_line22_FA2 ( l7_line22[3], l7_line22[4], l7_line22[5], l6_line22[6], l6_line23[1]) ;
   FA level7_line22_FA3 ( l7_line22[6], l7_line22[7], l7_line22[8], l6_line22[7], l6_line23[2]) ;
   FA level7_line22_FA4 ( l7_line22[9], l7_line22[10], l7_line22[11], l6_line22[8], l6_line23[3]) ;

   FA level7_line23_FA1 ( l7_line23[0], l7_line23[1], l7_line23[2], l6_line23[4], l6_line24[0]) ;
   FA level7_line23_FA2 ( l7_line23[3], l7_line23[4], l7_line23[5], l6_line23[5], l6_line24[1]) ;
   FA level7_line23_FA3 ( l7_line23[6], l7_line23[7], l7_line23[8], l6_line23[6], l6_line24[2]) ;

   FA level7_line24_FA1 ( l7_line24[0], l7_line24[1], l7_line24[2], l6_line24[3], l6_line25[0]) ;
   FA level7_line24_FA2 ( l7_line24[3], l7_line24[4], l7_line24[5], l6_line24[4], l6_line25[1]) ;

   FA level7_line25_FA1 ( l7_line25[0], l7_line25[1], l7_line25[2], l6_line25[2], l6_line26[0]) ;
	
	assign l6_line20[12] = l7_line20[17] ;
   assign l6_line21[12:11] = l7_line21[16:15] ;
   assign l6_line22[12:9] = l7_line22[15:12] ;
   assign l6_line23[12:7] = l7_line23[14:9] ;
   assign l6_line24[12:5] = l7_line24[13:6] ;
   assign l6_line25[12:3] = l7_line25[12:3] ;
	assign l6_line26[12:1] = l7_line26[11:0] ;
	
	// passing first 13 level 7 lines as it is to nect level with capacity of 13 wires
	assign l6_line1 = l7_line1 ;
   assign l6_line2 = l7_line2 ;
   assign l6_line3 = l7_line3 ;
   assign l6_line4 = l7_line4 ;
   assign l6_line5 = l7_line5 ;
   assign l6_line6 = l7_line6 ;
   assign l6_line7 = l7_line7 ;
   assign l6_line8 = l7_line8 ;
   assign l6_line9 = l7_line9 ;
   assign l6_line10 = l7_line10 ;
   assign l6_line11 = l7_line11 ;
   assign l6_line12 = l7_line12 ;
   assign l6_line13 = l7_line13 ;
	
	//passing rest of the values which will be passed to next level as it is
	assign l6_line27 = l7_line27 ;
   assign l6_line28 = l7_line28 ;
   assign l6_line29 = l7_line29 ;
   assign l6_line30 = l7_line30 ;
   assign l6_line31 = l7_line31 ;
   assign l6_line32 = l7_line32 ;
   assign l6_line33 = l7_line33 ;
   assign l6_line34 = l7_line34 ;
   assign l6_line35 = l7_line35 ;
   assign l6_line36 = l7_line36 ;
   assign l6_line37 = l7_line37 ;
	
	// Level-7 (19) to level-6 (13) complete
	// Declaring level-5 lines
	wire       l5_line1 ;
   wire [1:0] l5_line2 ;
   wire [2:0] l5_line3 ;
   wire [3:0] l5_line4 ;
   wire [4:0] l5_line5 ;
   wire [5:0] l5_line6 ;
   wire [6:0] l5_line7 ;
   wire [7:0] l5_line8 ;
   wire [8:0] l5_line9 ;
	
	wire [8:0] l5_line10 ;
   wire [8:0] l5_line11 ;
   wire [8:0] l5_line12 ;
   wire [8:0] l5_line13 ;
   wire [8:0] l5_line14 ;
   wire [8:0] l5_line15 ;
   wire [8:0] l5_line16 ;
   wire [8:0] l5_line17 ;
   wire [8:0] l5_line18 ;
   wire [8:0] l5_line19 ;
   wire [8:0] l5_line20 ;
   wire [8:0] l5_line21 ;
   wire [8:0] l5_line22 ;
   wire [8:0] l5_line23 ;
   wire [8:0] l5_line24 ;
   wire [8:0] l5_line25 ;
   wire [8:0] l5_line26 ;
   wire [8:0] l5_line27 ;
   wire [8:0] l5_line28 ;
   wire [8:0] l5_line29 ;
   wire [8:0] l5_line30 ;
	
	wire [6:0] l5_line31 ;
   wire [5:0] l5_line32 ;
   wire [4:0] l5_line33 ;
   wire [3:0] l5_line34 ;
   wire [2:0] l5_line35 ;
   wire [1:0] l5_line36 ;
   wire [0:0] l5_line37 ;
	
	// instantiating ful adders for level-5 in level-6
	HA level6_line10_HA1 ( l6_line10[0], l6_line10[1],              l5_line10[0], l5_line11[0]) ;
	
   FA level6_line11_FA1 ( l6_line11[0], l6_line11[1], l6_line11[2], l5_line11[1], l5_line12[0]) ;
   HA level6_line11_HA1 ( l6_line11[3], l6_line11[4],              l5_line11[2], l5_line12[1]) ;

   FA level6_line12_FA1 ( l6_line12[0], l6_line12[1], l6_line12[2], l5_line12[2], l5_line13[0]) ;
   FA level6_line12_FA2 ( l6_line12[3], l6_line12[4], l6_line12[5], l5_line12[3], l5_line13[1]) ;
   HA level6_line12_HA1 ( l6_line12[6], l6_line12[7],              l5_line12[4], l5_line13[2]) ;

   FA level6_line13_FA1 ( l6_line13[0], l6_line13[1], l6_line13[2], l5_line13[3], l5_line14[0]) ;
   FA level6_line13_FA2 ( l6_line13[3], l6_line13[4], l6_line13[5], l5_line13[4], l5_line14[1]) ;
   FA level6_line13_FA3 ( l6_line13[6], l6_line13[7], l6_line13[8], l5_line13[5], l5_line14[2]) ;
   HA level6_line13_HA1 ( l6_line13[9], l6_line13[10],              l5_line13[6], l5_line14[3]) ;
	
	assign l5_line10[8:1] = l6_line10[9:2] ;
   assign l5_line11[8:3] = l6_line11[10:5] ;
   assign l5_line12[8:5] = l6_line12[11:8] ;
   assign l5_line13[8:7] = l6_line13[12:11] ;
	
   FA level6_line14_FA1 ( l6_line14[0], l6_line14[1], l6_line14[2], l5_line14[4], l5_line15[0]) ;
   FA level6_line14_FA2 ( l6_line14[3], l6_line14[4], l6_line14[5], l5_line14[5], l5_line15[1]) ;
   FA level6_line14_FA3 ( l6_line14[6], l6_line14[7], l6_line14[8], l5_line14[6], l5_line15[2]) ;
   FA level6_line14_FA4 ( l6_line14[9], l6_line14[10], l6_line14[11], l5_line14[7], l5_line15[3]) ;

   FA level6_line15_FA1 ( l6_line15[0], l6_line15[1], l6_line15[2], l5_line15[4], l5_line16[0]) ;
   FA level6_line15_FA2 ( l6_line15[3], l6_line15[4], l6_line15[5], l5_line15[5], l5_line16[1]) ;
   FA level6_line15_FA3 ( l6_line15[6], l6_line15[7], l6_line15[8], l5_line15[6], l5_line16[2]) ;
   FA level6_line15_FA4 ( l6_line15[9], l6_line15[10], l6_line15[11], l5_line15[7], l5_line16[3]) ;

   FA level6_line16_FA1 ( l6_line16[0], l6_line16[1], l6_line16[2], l5_line16[4], l5_line17[0]) ;
   FA level6_line16_FA2 ( l6_line16[3], l6_line16[4], l6_line16[5], l5_line16[5], l5_line17[1]) ;
   FA level6_line16_FA3 ( l6_line16[6], l6_line16[7], l6_line16[8], l5_line16[6], l5_line17[2]) ;
   FA level6_line16_FA4 ( l6_line16[9], l6_line16[10], l6_line16[11], l5_line16[7], l5_line17[3]) ;

   FA level6_line17_FA1 ( l6_line17[0], l6_line17[1], l6_line17[2], l5_line17[4], l5_line18[0]) ;
   FA level6_line17_FA2 ( l6_line17[3], l6_line17[4], l6_line17[5], l5_line17[5], l5_line18[1]) ;
   FA level6_line17_FA3 ( l6_line17[6], l6_line17[7], l6_line17[8], l5_line17[6], l5_line18[2]) ;
   FA level6_line17_FA4 ( l6_line17[9], l6_line17[10], l6_line17[11], l5_line17[7], l5_line18[3]) ;

   FA level6_line18_FA1 ( l6_line18[0], l6_line18[1], l6_line18[2], l5_line18[4], l5_line19[0]) ;
   FA level6_line18_FA2 ( l6_line18[3], l6_line18[4], l6_line18[5], l5_line18[5], l5_line19[1]) ;
   FA level6_line18_FA3 ( l6_line18[6], l6_line18[7], l6_line18[8], l5_line18[6], l5_line19[2]) ;
   FA level6_line18_FA4 ( l6_line18[9], l6_line18[10], l6_line18[11], l5_line18[7], l5_line19[3]) ;

   FA level6_line19_FA1 ( l6_line19[0], l6_line19[1], l6_line19[2], l5_line19[4], l5_line20[0]) ;
   FA level6_line19_FA2 ( l6_line19[3], l6_line19[4], l6_line19[5], l5_line19[5], l5_line20[1]) ;
   FA level6_line19_FA3 ( l6_line19[6], l6_line19[7], l6_line19[8], l5_line19[6], l5_line20[2]) ;
   FA level6_line19_FA4 ( l6_line19[9], l6_line19[10], l6_line19[11], l5_line19[7], l5_line20[3]) ;

   FA level6_line20_FA1 ( l6_line20[0], l6_line20[1], l6_line20[2], l5_line20[4], l5_line21[0]) ;
   FA level6_line20_FA2 ( l6_line20[3], l6_line20[4], l6_line20[5], l5_line20[5], l5_line21[1]) ;
   FA level6_line20_FA3 ( l6_line20[6], l6_line20[7], l6_line20[8], l5_line20[6], l5_line21[2]) ;
   FA level6_line20_FA4 ( l6_line20[9], l6_line20[10], l6_line20[11], l5_line20[7], l5_line21[3]) ;

   FA level6_line21_FA1 ( l6_line21[0], l6_line21[1], l6_line21[2], l5_line21[4], l5_line22[0]) ;
   FA level6_line21_FA2 ( l6_line21[3], l6_line21[4], l6_line21[5], l5_line21[5], l5_line22[1]) ;
   FA level6_line21_FA3 ( l6_line21[6], l6_line21[7], l6_line21[8], l5_line21[6], l5_line22[2]) ;
   FA level6_line21_FA4 ( l6_line21[9], l6_line21[10], l6_line21[11], l5_line21[7], l5_line22[3]) ;

   FA level6_line22_FA1 ( l6_line22[0], l6_line22[1], l6_line22[2], l5_line22[4], l5_line23[0]) ;
   FA level6_line22_FA2 ( l6_line22[3], l6_line22[4], l6_line22[5], l5_line22[5], l5_line23[1]) ;
   FA level6_line22_FA3 ( l6_line22[6], l6_line22[7], l6_line22[8], l5_line22[6], l5_line23[2]) ;
   FA level6_line22_FA4 ( l6_line22[9], l6_line22[10], l6_line22[11], l5_line22[7], l5_line23[3]) ;

   FA level6_line23_FA1 ( l6_line23[0], l6_line23[1], l6_line23[2], l5_line23[4], l5_line24[0]) ;
   FA level6_line23_FA2 ( l6_line23[3], l6_line23[4], l6_line23[5], l5_line23[5], l5_line24[1]) ;
   FA level6_line23_FA3 ( l6_line23[6], l6_line23[7], l6_line23[8], l5_line23[6], l5_line24[2]) ;
   FA level6_line23_FA4 ( l6_line23[9], l6_line23[10], l6_line23[11], l5_line23[7], l5_line24[3]) ;

   FA level6_line24_FA1 ( l6_line24[0], l6_line24[1], l6_line24[2], l5_line24[4], l5_line25[0]) ;
   FA level6_line24_FA2 ( l6_line24[3], l6_line24[4], l6_line24[5], l5_line24[5], l5_line25[1]) ;
   FA level6_line24_FA3 ( l6_line24[6], l6_line24[7], l6_line24[8], l5_line24[6], l5_line25[2]) ;
   FA level6_line24_FA4 ( l6_line24[9], l6_line24[10], l6_line24[11], l5_line24[7], l5_line25[3]) ;

   FA level6_line25_FA1 ( l6_line25[0], l6_line25[1], l6_line25[2], l5_line25[4], l5_line26[0]) ;
   FA level6_line25_FA2 ( l6_line25[3], l6_line25[4], l6_line25[5], l5_line25[5], l5_line26[1]) ;
   FA level6_line25_FA3 ( l6_line25[6], l6_line25[7], l6_line25[8], l5_line25[6], l5_line26[2]) ;
   FA level6_line25_FA4 ( l6_line25[9], l6_line25[10], l6_line25[11], l5_line25[7], l5_line26[3]) ;
	
   FA level6_line26_FA1 ( l6_line26[0], l6_line26[1], l6_line26[2], l5_line26[4], l5_line27[0]) ;
   FA level6_line26_FA2 ( l6_line26[3], l6_line26[4], l6_line26[5], l5_line26[5], l5_line27[1]) ;
   FA level6_line26_FA3 ( l6_line26[6], l6_line26[7], l6_line26[8], l5_line26[6], l5_line27[2]) ;
   FA level6_line26_FA4 ( l6_line26[9], l6_line26[10], l6_line26[11], l5_line26[7], l5_line27[3]) ;
	
	assign l5_line14[8] = l6_line14[12] ;
   assign l5_line15[8] = l6_line15[12] ;
   assign l5_line16[8] = l6_line16[12] ;
   assign l5_line17[8] = l6_line17[12] ;
   assign l5_line18[8] = l6_line18[12] ;
   assign l5_line19[8] = l6_line19[12] ;
   assign l5_line20[8] = l6_line20[12] ;
   assign l5_line21[8] = l6_line21[12] ;
   assign l5_line22[8] = l6_line22[12] ;
   assign l5_line23[8] = l6_line23[12] ;
   assign l5_line24[8] = l6_line24[12] ;
   assign l5_line25[8] = l6_line25[12] ;
   assign l5_line26[8] = l6_line26[12] ;
	
   FA level6_line27_FA1 ( l6_line27[0], l6_line27[1], l6_line27[2], l5_line27[4], l5_line28[0]) ;
   FA level6_line27_FA2 ( l6_line27[3], l6_line27[4], l6_line27[5], l5_line27[5], l5_line28[1]) ;
   FA level6_line27_FA3 ( l6_line27[6], l6_line27[7], l6_line27[8], l5_line27[6], l5_line28[2]) ;

   FA level6_line28_FA1 ( l6_line28[0], l6_line28[1], l6_line28[2], l5_line28[3], l5_line29[0]) ;
   FA level6_line28_FA2 ( l6_line28[3], l6_line28[4], l6_line28[5], l5_line28[4], l5_line29[1]) ;

   FA level6_line29_FA1 ( l6_line29[0], l6_line29[1], l6_line29[2], l5_line29[2], l5_line30[0]) ;
	
	assign l5_line27[8:7] = l6_line27[10:9] ;
   assign l5_line28[8:5] = l6_line28[9:6] ;
   assign l5_line29[8:3] = l6_line29[8:3] ;
   assign l5_line30[8:1] = l6_line30[7:0] ;
	
	// passing first 13 level 7 lines as it is to nect level with capacity of 13 wires
	assign l5_line1 = l6_line1 ;
   assign l5_line2 = l6_line2 ;
   assign l5_line3 = l6_line3 ;
   assign l5_line4 = l6_line4 ;
   assign l5_line5 = l6_line5 ;
   assign l5_line6 = l6_line6 ;
   assign l5_line7 = l6_line7 ;
   assign l5_line8 = l6_line8 ;
   assign l5_line9 = l6_line9 ;
	
	//passing rest of the values which will be passed to next level as it is
   assign l5_line31 = l6_line31 ;
   assign l5_line32 = l6_line32 ;
   assign l5_line33 = l6_line33 ;
   assign l5_line34 = l6_line34 ;
   assign l5_line35 = l6_line35 ;
   assign l5_line36 = l6_line36 ;
   assign l5_line37 = l6_line37 ;
	
	// Level-6 (13) to level-5 (9) complete
	// Declaring level-4 lines
	wire       l4_line1 ;
   wire [1:0] l4_line2 ;
   wire [2:0] l4_line3 ;
   wire [3:0] l4_line4 ;
   wire [4:0] l4_line5 ;
   wire [5:0] l4_line6 ;
	
   wire [5:0] l4_line7 ;
   wire [5:0] l4_line8 ;
   wire [5:0] l4_line9 ;
   wire [5:0] l4_line10 ;
   wire [5:0] l4_line11 ;
   wire [5:0] l4_line12 ;
   wire [5:0] l4_line13 ;
   wire [5:0] l4_line14 ;
   wire [5:0] l4_line15 ;
   wire [5:0] l4_line16 ;
   wire [5:0] l4_line17 ;
   wire [5:0] l4_line18 ;
   wire [5:0] l4_line19 ;
   wire [5:0] l4_line20 ;
   wire [5:0] l4_line21 ;
   wire [5:0] l4_line22 ;
   wire [5:0] l4_line23 ;
   wire [5:0] l4_line24 ;
   wire [5:0] l4_line25 ;
   wire [5:0] l4_line26 ;
   wire [5:0] l4_line27 ;
   wire [5:0] l4_line28 ;
   wire [5:0] l4_line29 ;
   wire [5:0] l4_line30 ;
   wire [5:0] l4_line31 ;
   wire [5:0] l4_line32 ;
   wire [5:0] l4_line33 ;
	
   wire [3:0] l4_line34 ;
   wire [2:0] l4_line35 ;
   wire [1:0] l4_line36 ;
   wire       l4_line37 ;
	
	// instantiating ful adders for level-4 in level-5
	HA level5_line7_HA1 ( l5_line7[0], l5_line7[1],              l4_line7[0], l4_line8[0]) ;

   FA level5_line8_FA1 ( l5_line8[0], l5_line8[1], l5_line8[2], l4_line8[1], l4_line9[0]) ;
   HA level5_line8_HA1 ( l5_line8[3], l5_line8[4],              l4_line8[2], l4_line9[1]) ;

   FA level5_line9_FA1 ( l5_line9[0], l5_line9[1], l5_line9[2], l4_line9[2], l4_line10[0]) ;
   FA level5_line9_FA2 ( l5_line9[3], l5_line9[4], l5_line9[5], l4_line9[3], l4_line10[1]) ;
   HA level5_line9_HA1 ( l5_line9[6], l5_line9[7],              l4_line9[4], l4_line10[2]) ;
	
	assign l4_line7[5:1] = l5_line7[6:2] ;
   assign l4_line8[5:3] = l5_line8[7:5] ;
   assign l4_line9[5] = l5_line9[8] ;
	
   FA level5_line10_FA1 ( l5_line10[0], l5_line10[1], l5_line10[2], l4_line10[3], l4_line11[0]) ;
   FA level5_line10_FA2 ( l5_line10[3], l5_line10[4], l5_line10[5], l4_line10[4], l4_line11[1]) ;
   FA level5_line10_FA3 ( l5_line10[6], l5_line10[7], l5_line10[8], l4_line10[5], l4_line11[2]) ;

   FA level5_line11_FA1 ( l5_line11[0], l5_line11[1], l5_line11[2], l4_line11[3], l4_line12[0]) ;
   FA level5_line11_FA2 ( l5_line11[3], l5_line11[4], l5_line11[5], l4_line11[4], l4_line12[1]) ;
   FA level5_line11_FA3 ( l5_line11[6], l5_line11[7], l5_line11[8], l4_line11[5], l4_line12[2]) ;

   FA level5_line12_FA1 ( l5_line12[0], l5_line12[1], l5_line12[2], l4_line12[3], l4_line13[0]) ;
   FA level5_line12_FA2 ( l5_line12[3], l5_line12[4], l5_line12[5], l4_line12[4], l4_line13[1]) ;
   FA level5_line12_FA3 ( l5_line12[6], l5_line12[7], l5_line12[8], l4_line12[5], l4_line13[2]) ;

   FA level5_line13_FA1 ( l5_line13[0], l5_line13[1], l5_line13[2], l4_line13[3], l4_line14[0]) ;
   FA level5_line13_FA2 ( l5_line13[3], l5_line13[4], l5_line13[5], l4_line13[4], l4_line14[1]) ;
   FA level5_line13_FA3 ( l5_line13[6], l5_line13[7], l5_line13[8], l4_line13[5], l4_line14[2]) ;

   FA level5_line14_FA1 ( l5_line14[0], l5_line14[1], l5_line14[2], l4_line14[3], l4_line15[0]) ;
   FA level5_line14_FA2 ( l5_line14[3], l5_line14[4], l5_line14[5], l4_line14[4], l4_line15[1]) ;
   FA level5_line14_FA3 ( l5_line14[6], l5_line14[7], l5_line14[8], l4_line14[5], l4_line15[2]) ;

   FA level5_line15_FA1 ( l5_line15[0], l5_line15[1], l5_line15[2], l4_line15[3], l4_line16[0]) ;
   FA level5_line15_FA2 ( l5_line15[3], l5_line15[4], l5_line15[5], l4_line15[4], l4_line16[1]) ;
   FA level5_line15_FA3 ( l5_line15[6], l5_line15[7], l5_line15[8], l4_line15[5], l4_line16[2]) ;

   FA level5_line16_FA1 ( l5_line16[0], l5_line16[1], l5_line16[2], l4_line16[3], l4_line17[0]) ;
   FA level5_line16_FA2 ( l5_line16[3], l5_line16[4], l5_line16[5], l4_line16[4], l4_line17[1]) ;
   FA level5_line16_FA3 ( l5_line16[6], l5_line16[7], l5_line16[8], l4_line16[5], l4_line17[2]) ;

   FA level5_line17_FA1 ( l5_line17[0], l5_line17[1], l5_line17[2], l4_line17[3], l4_line18[0]) ;
   FA level5_line17_FA2 ( l5_line17[3], l5_line17[4], l5_line17[5], l4_line17[4], l4_line18[1]) ;
   FA level5_line17_FA3 ( l5_line17[6], l5_line17[7], l5_line17[8], l4_line17[5], l4_line18[2]) ;

   FA level5_line18_FA1 ( l5_line18[0], l5_line18[1], l5_line18[2], l4_line18[3], l4_line19[0]) ;
   FA level5_line18_FA2 ( l5_line18[3], l5_line18[4], l5_line18[5], l4_line18[4], l4_line19[1]) ;
   FA level5_line18_FA3 ( l5_line18[6], l5_line18[7], l5_line18[8], l4_line18[5], l4_line19[2]) ;

   FA level5_line19_FA1 ( l5_line19[0], l5_line19[1], l5_line19[2], l4_line19[3], l4_line20[0]) ;
   FA level5_line19_FA2 ( l5_line19[3], l5_line19[4], l5_line19[5], l4_line19[4], l4_line20[1]) ;
   FA level5_line19_FA3 ( l5_line19[6], l5_line19[7], l5_line19[8], l4_line19[5], l4_line20[2]) ;

   FA level5_line20_FA1 ( l5_line20[0], l5_line20[1], l5_line20[2], l4_line20[3], l4_line21[0]) ;
   FA level5_line20_FA2 ( l5_line20[3], l5_line20[4], l5_line20[5], l4_line20[4], l4_line21[1]) ;
   FA level5_line20_FA3 ( l5_line20[6], l5_line20[7], l5_line20[8], l4_line20[5], l4_line21[2]) ;

   FA level5_line21_FA1 ( l5_line21[0], l5_line21[1], l5_line21[2], l4_line21[3], l4_line22[0]) ;
   FA level5_line21_FA2 ( l5_line21[3], l5_line21[4], l5_line21[5], l4_line21[4], l4_line22[1]) ;
   FA level5_line21_FA3 ( l5_line21[6], l5_line21[7], l5_line21[8], l4_line21[5], l4_line22[2]) ;

   FA level5_line22_FA1 ( l5_line22[0], l5_line22[1], l5_line22[2], l4_line22[3], l4_line23[0]) ;
   FA level5_line22_FA2 ( l5_line22[3], l5_line22[4], l5_line22[5], l4_line22[4], l4_line23[1]) ;
   FA level5_line22_FA3 ( l5_line22[6], l5_line22[7], l5_line22[8], l4_line22[5], l4_line23[2]) ;

   FA level5_line23_FA1 ( l5_line23[0], l5_line23[1], l5_line23[2], l4_line23[3], l4_line24[0]) ;
   FA level5_line23_FA2 ( l5_line23[3], l5_line23[4], l5_line23[5], l4_line23[4], l4_line24[1]) ;
   FA level5_line23_FA3 ( l5_line23[6], l5_line23[7], l5_line23[8], l4_line23[5], l4_line24[2]) ;

   FA level5_line24_FA1 ( l5_line24[0], l5_line24[1], l5_line24[2], l4_line24[3], l4_line25[0]) ;
   FA level5_line24_FA2 ( l5_line24[3], l5_line24[4], l5_line24[5], l4_line24[4], l4_line25[1]) ;
   FA level5_line24_FA3 ( l5_line24[6], l5_line24[7], l5_line24[8], l4_line24[5], l4_line25[2]) ;

   FA level5_line25_FA1 ( l5_line25[0], l5_line25[1], l5_line25[2], l4_line25[3], l4_line26[0]) ;
   FA level5_line25_FA2 ( l5_line25[3], l5_line25[4], l5_line25[5], l4_line25[4], l4_line26[1]) ;
   FA level5_line25_FA3 ( l5_line25[6], l5_line25[7], l5_line25[8], l4_line25[5], l4_line26[2]) ;

   FA level5_line26_FA1 ( l5_line26[0], l5_line26[1], l5_line26[2], l4_line26[3], l4_line27[0]) ;
   FA level5_line26_FA2 ( l5_line26[3], l5_line26[4], l5_line26[5], l4_line26[4], l4_line27[1]) ;
   FA level5_line26_FA3 ( l5_line26[6], l5_line26[7], l5_line26[8], l4_line26[5], l4_line27[2]) ;

   FA level5_line27_FA1 ( l5_line27[0], l5_line27[1], l5_line27[2], l4_line27[3], l4_line28[0]) ;
   FA level5_line27_FA2 ( l5_line27[3], l5_line27[4], l5_line27[5], l4_line27[4], l4_line28[1]) ;
   FA level5_line27_FA3 ( l5_line27[6], l5_line27[7], l5_line27[8], l4_line27[5], l4_line28[2]) ;

   FA level5_line28_FA1 ( l5_line28[0], l5_line28[1], l5_line28[2], l4_line28[3], l4_line29[0]) ;
   FA level5_line28_FA2 ( l5_line28[3], l5_line28[4], l5_line28[5], l4_line28[4], l4_line29[1]) ;
   FA level5_line28_FA3 ( l5_line28[6], l5_line28[7], l5_line28[8], l4_line28[5], l4_line29[2]) ;

   FA level5_line29_FA1 ( l5_line29[0], l5_line29[1], l5_line29[2], l4_line29[3], l4_line30[0]) ;
   FA level5_line29_FA2 ( l5_line29[3], l5_line29[4], l5_line29[5], l4_line29[4], l4_line30[1]) ;
   FA level5_line29_FA3 ( l5_line29[6], l5_line29[7], l5_line29[8], l4_line29[5], l4_line30[2]) ;

   FA level5_line30_FA1 ( l5_line30[0], l5_line30[1], l5_line30[2], l4_line30[3], l4_line31[0]) ;
   FA level5_line30_FA2 ( l5_line30[3], l5_line30[4], l5_line30[5], l4_line30[4], l4_line31[1]) ;
   FA level5_line30_FA3 ( l5_line30[6], l5_line30[7], l5_line30[8], l4_line30[5], l4_line31[2]) ;

   FA level5_line31_FA1 ( l5_line31[0], l5_line31[1], l5_line31[2], l4_line31[3], l4_line32[0]) ;
   FA level5_line31_FA2 ( l5_line31[3], l5_line31[4], l5_line31[5], l4_line31[4], l4_line32[1]) ;

   FA level5_line32_FA1 ( l5_line32[0], l5_line32[1], l5_line32[2], l4_line32[2], l4_line33[0]) ;
	
	assign l4_line31[5] = l5_line31[6] ;
	assign l4_line32[5:3] = l5_line32[5:3] ;
	assign l4_line33[5:1] = l5_line33[4:0] ;
	
	// passing first 6 level 5 lines as it is to nect level with capacity of 6 wires
	assign l4_line1 = l5_line1 ;
   assign l4_line2 = l5_line2 ;
   assign l4_line3 = l5_line3 ;
   assign l4_line4 = l5_line4 ;
   assign l4_line5 = l5_line5 ;
   assign l4_line6 = l5_line6 ;
	
	//passing rest of the values which will be passed to next level as it is
   assign l4_line34 = l5_line34 ;
   assign l4_line35 = l5_line35 ;
   assign l4_line36 = l5_line36 ;
   assign l4_line37 = l5_line37 ;
	
	// Level-5 (9) to level-4 (6) complete
	// Declaring level-3 lines
	wire 	     l3_line1 ;
   wire [1:0] l3_line2 ;
   wire [2:0] l3_line3 ;
   wire [3:0] l3_line4 ;
	
   wire [3:0] l3_line5 ;
   wire [3:0] l3_line6 ;
   wire [3:0] l3_line7 ;
   wire [3:0] l3_line8 ;
   wire [3:0] l3_line9 ;
   wire [3:0] l3_line10 ;
   wire [3:0] l3_line11 ;
   wire [3:0] l3_line12 ;
   wire [3:0] l3_line13 ;
   wire [3:0] l3_line14 ;
   wire [3:0] l3_line15 ;
   wire [3:0] l3_line16 ;
   wire [3:0] l3_line17 ;
   wire [3:0] l3_line18 ;
   wire [3:0] l3_line19 ;
   wire [3:0] l3_line20 ;
   wire [3:0] l3_line21 ;
   wire [3:0] l3_line22 ;
   wire [3:0] l3_line23 ;
   wire [3:0] l3_line24 ;
   wire [3:0] l3_line25 ;
   wire [3:0] l3_line26 ;
   wire [3:0] l3_line27 ;
   wire [3:0] l3_line28 ;
   wire [3:0] l3_line29 ;
   wire [3:0] l3_line30 ;
   wire [3:0] l3_line31 ;
   wire [3:0] l3_line32 ;
   wire [3:0] l3_line33 ;
   wire [3:0] l3_line34 ;
   wire [3:0] l3_line35 ;
	
   wire [1:0] l3_line36 ;
   wire       l3_line37 ;
	
	// instantiating ful adders for level-3 in level-4
	HA level4_line5_HA1 ( l4_line5[0], l4_line5[1],              l3_line5[0], l3_line6[0]) ;
	
   FA level4_line6_FA1 ( l4_line6[0], l4_line6[1], l4_line6[2], l3_line6[1], l3_line7[0]) ;
   HA level4_line6_HA1 ( l4_line6[3], l4_line6[4],              l3_line6[2], l3_line7[1]) ;

   FA level4_line7_FA1 ( l4_line7[0], l4_line7[1], l4_line7[2], l3_line7[2], l3_line8[0]) ;
   FA level4_line7_FA2 ( l4_line7[3], l4_line7[4], l4_line7[5], l3_line7[3], l3_line8[1]) ;

   FA level4_line8_FA1 ( l4_line8[0], l4_line8[1], l4_line8[2], l3_line8[2], l3_line9[0]) ;
   FA level4_line8_FA2 ( l4_line8[3], l4_line8[4], l4_line8[5], l3_line8[3], l3_line9[1]) ;

   FA level4_line9_FA1 ( l4_line9[0], l4_line9[1], l4_line9[2], l3_line9[2], l3_line10[0]) ;
   FA level4_line9_FA2 ( l4_line9[3], l4_line9[4], l4_line9[5], l3_line9[3], l3_line10[1]) ;

   FA level4_line10_FA1 ( l4_line10[0], l4_line10[1], l4_line10[2], l3_line10[2], l3_line11[0]) ;
   FA level4_line10_FA2 ( l4_line10[3], l4_line10[4], l4_line10[5], l3_line10[3], l3_line11[1]) ;

   FA level4_line11_FA1 ( l4_line11[0], l4_line11[1], l4_line11[2], l3_line11[2], l3_line12[0]) ;
   FA level4_line11_FA2 ( l4_line11[3], l4_line11[4], l4_line11[5], l3_line11[3], l3_line12[1]) ;

   FA level4_line12_FA1 ( l4_line12[0], l4_line12[1], l4_line12[2], l3_line12[2], l3_line13[0]) ;
   FA level4_line12_FA2 ( l4_line12[3], l4_line12[4], l4_line12[5], l3_line12[3], l3_line13[1]) ;

   FA level4_line13_FA1 ( l4_line13[0], l4_line13[1], l4_line13[2], l3_line13[2], l3_line14[0]) ;
   FA level4_line13_FA2 ( l4_line13[3], l4_line13[4], l4_line13[5], l3_line13[3], l3_line14[1]) ;

   FA level4_line14_FA1 ( l4_line14[0], l4_line14[1], l4_line14[2], l3_line14[2], l3_line15[0]) ;
   FA level4_line14_FA2 ( l4_line14[3], l4_line14[4], l4_line14[5], l3_line14[3], l3_line15[1]) ;

   FA level4_line15_FA1 ( l4_line15[0], l4_line15[1], l4_line15[2], l3_line15[2], l3_line16[0]) ;
   FA level4_line15_FA2 ( l4_line15[3], l4_line15[4], l4_line15[5], l3_line15[3], l3_line16[1]) ;

   FA level4_line16_FA1 ( l4_line16[0], l4_line16[1], l4_line16[2], l3_line16[2], l3_line17[0]) ;
   FA level4_line16_FA2 ( l4_line16[3], l4_line16[4], l4_line16[5], l3_line16[3], l3_line17[1]) ;

   FA level4_line17_FA1 ( l4_line17[0], l4_line17[1], l4_line17[2], l3_line17[2], l3_line18[0]) ;
   FA level4_line17_FA2 ( l4_line17[3], l4_line17[4], l4_line17[5], l3_line17[3], l3_line18[1]) ;

   FA level4_line18_FA1 ( l4_line18[0], l4_line18[1], l4_line18[2], l3_line18[2], l3_line19[0]) ;
   FA level4_line18_FA2 ( l4_line18[3], l4_line18[4], l4_line18[5], l3_line18[3], l3_line19[1]) ;

   FA level4_line19_FA1 ( l4_line19[0], l4_line19[1], l4_line19[2], l3_line19[2], l3_line20[0]) ;
   FA level4_line19_FA2 ( l4_line19[3], l4_line19[4], l4_line19[5], l3_line19[3], l3_line20[1]) ;

   FA level4_line20_FA1 ( l4_line20[0], l4_line20[1], l4_line20[2], l3_line20[2], l3_line21[0]) ;
   FA level4_line20_FA2 ( l4_line20[3], l4_line20[4], l4_line20[5], l3_line20[3], l3_line21[1]) ;

   FA level4_line21_FA1 ( l4_line21[0], l4_line21[1], l4_line21[2], l3_line21[2], l3_line22[0]) ;
   FA level4_line21_FA2 ( l4_line21[3], l4_line21[4], l4_line21[5], l3_line21[3], l3_line22[1]) ;

   FA level4_line22_FA1 ( l4_line22[0], l4_line22[1], l4_line22[2], l3_line22[2], l3_line23[0]) ;
   FA level4_line22_FA2 ( l4_line22[3], l4_line22[4], l4_line22[5], l3_line22[3], l3_line23[1]) ;

   FA level4_line23_FA1 ( l4_line23[0], l4_line23[1], l4_line23[2], l3_line23[2], l3_line24[0]) ;
   FA level4_line23_FA2 ( l4_line23[3], l4_line23[4], l4_line23[5], l3_line23[3], l3_line24[1]) ;

   FA level4_line24_FA1 ( l4_line24[0], l4_line24[1], l4_line24[2], l3_line24[2], l3_line25[0]) ;
   FA level4_line24_FA2 ( l4_line24[3], l4_line24[4], l4_line24[5], l3_line24[3], l3_line25[1]) ;

   FA level4_line25_FA1 ( l4_line25[0], l4_line25[1], l4_line25[2], l3_line25[2], l3_line26[0]) ;
   FA level4_line25_FA2 ( l4_line25[3], l4_line25[4], l4_line25[5], l3_line25[3], l3_line26[1]) ;

   FA level4_line26_FA1 ( l4_line26[0], l4_line26[1], l4_line26[2], l3_line26[2], l3_line27[0]) ;
   FA level4_line26_FA2 ( l4_line26[3], l4_line26[4], l4_line26[5], l3_line26[3], l3_line27[1]) ;

   FA level4_line27_FA1 ( l4_line27[0], l4_line27[1], l4_line27[2], l3_line27[2], l3_line28[0]) ;
   FA level4_line27_FA2 ( l4_line27[3], l4_line27[4], l4_line27[5], l3_line27[3], l3_line28[1]) ;

   FA level4_line28_FA1 ( l4_line28[0], l4_line28[1], l4_line28[2], l3_line28[2], l3_line29[0]) ;
   FA level4_line28_FA2 ( l4_line28[3], l4_line28[4], l4_line28[5], l3_line28[3], l3_line29[1]) ;

   FA level4_line29_FA1 ( l4_line29[0], l4_line29[1], l4_line29[2], l3_line29[2], l3_line30[0]) ;
   FA level4_line29_FA2 ( l4_line29[3], l4_line29[4], l4_line29[5], l3_line29[3], l3_line30[1]) ;

   FA level4_line30_FA1 ( l4_line30[0], l4_line30[1], l4_line30[2], l3_line30[2], l3_line31[0]) ;
   FA level4_line30_FA2 ( l4_line30[3], l4_line30[4], l4_line30[5], l3_line30[3], l3_line31[1]) ;

   FA level4_line31_FA1 ( l4_line31[0], l4_line31[1], l4_line31[2], l3_line31[2], l3_line32[0]) ;
   FA level4_line31_FA2 ( l4_line31[3], l4_line31[4], l4_line31[5], l3_line31[3], l3_line32[1]) ;

   FA level4_line32_FA1 ( l4_line32[0], l4_line32[1], l4_line32[2], l3_line32[2], l3_line33[0]) ;
   FA level4_line32_FA2 ( l4_line32[3], l4_line32[4], l4_line32[5], l3_line32[3], l3_line33[1]) ;

   FA level4_line33_FA1 ( l4_line33[0], l4_line33[1], l4_line33[2], l3_line33[2], l3_line34[0]) ;
   FA level4_line33_FA2 ( l4_line33[3], l4_line33[4], l4_line33[5], l3_line33[3], l3_line34[1]) ;

   FA level4_line34_FA1 ( l4_line34[0], l4_line34[1], l4_line34[2], l3_line34[2], l3_line35[0]) ;
	
	assign l3_line5[3:1] = l4_line5[4:2] ;
   assign l3_line6[3] = l4_line6[5] ;
	
	assign l3_line34[3] = l4_line34[3] ;
	assign l3_line35[3:1] = l4_line35[2:0] ;
	
	// passing first 4 level 4 lines as it is to nect level with capacity of 4 wires
	assign l3_line1 = l4_line1 ;
   assign l3_line2 = l4_line2 ;
   assign l3_line3 = l4_line3 ;
   assign l3_line4 = l4_line4 ;
	
	//passing rest of the values which will be passed to next level as it is
   assign l3_line36 = l4_line36 ;
   assign l3_line37 = l4_line37 ;
	
	// Level-4 (6) to level-3 (4) complete
	// Declaring level-2 lines
	wire       l2_line1 ;
   wire [1:0] l2_line2 ;
   wire [2:0] l2_line3 ;
	
   wire [2:0] l2_line4 ;
   wire [2:0] l2_line5 ;
   wire [2:0] l2_line6 ;
   wire [2:0] l2_line7 ;
   wire [2:0] l2_line8 ;
   wire [2:0] l2_line9 ;
   wire [2:0] l2_line10 ;
   wire [2:0] l2_line11 ;
   wire [2:0] l2_line12 ;
   wire [2:0] l2_line13 ;
   wire [2:0] l2_line14 ;
   wire [2:0] l2_line15 ;
   wire [2:0] l2_line16 ;
   wire [2:0] l2_line17 ;
   wire [2:0] l2_line18 ;
   wire [2:0] l2_line19 ;
   wire [2:0] l2_line20 ;
   wire [2:0] l2_line21 ;
   wire [2:0] l2_line22 ;
   wire [2:0] l2_line23 ;
   wire [2:0] l2_line24 ;
   wire [2:0] l2_line25 ;
   wire [2:0] l2_line26 ;
   wire [2:0] l2_line27 ;
   wire [2:0] l2_line28 ;
   wire [2:0] l2_line29 ;
   wire [2:0] l2_line30 ;
   wire [2:0] l2_line31 ;
   wire [2:0] l2_line32 ;
   wire [2:0] l2_line33 ;
   wire [2:0] l2_line34 ;
   wire [2:0] l2_line35 ;
   wire [2:0] l2_line36 ;
	
   wire       l2_line37 ;
	
	// instantiating ful adders for level-3 in level-4
	HA level3_line4_HA1 ( l3_line4[0], l3_line4[1],              l2_line4[0], l2_line5[0]) ;
	assign l2_line4[2:1] = l3_line4[3:2] ;
	
   FA level3_line5_FA1 ( l3_line5[0], l3_line5[1], l3_line5[2], l2_line5[1], l2_line6[0]) ;

   FA level3_line6_FA1 ( l3_line6[0], l3_line6[1], l3_line6[2], l2_line6[1], l2_line7[0]) ;

   FA level3_line7_FA1 ( l3_line7[0], l3_line7[1], l3_line7[2], l2_line7[1], l2_line8[0]) ;

   FA level3_line8_FA1 ( l3_line8[0], l3_line8[1], l3_line8[2], l2_line8[1], l2_line9[0]) ;

   FA level3_line9_FA1 ( l3_line9[0], l3_line9[1], l3_line9[2], l2_line9[1], l2_line10[0]) ;

   FA level3_line10_FA1 ( l3_line10[0], l3_line10[1], l3_line10[2], l2_line10[1], l2_line11[0]) ;

   FA level3_line11_FA1 ( l3_line11[0], l3_line11[1], l3_line11[2], l2_line11[1], l2_line12[0]) ;

   FA level3_line12_FA1 ( l3_line12[0], l3_line12[1], l3_line12[2], l2_line12[1], l2_line13[0]) ;

   FA level3_line13_FA1 ( l3_line13[0], l3_line13[1], l3_line13[2], l2_line13[1], l2_line14[0]) ;

   FA level3_line14_FA1 ( l3_line14[0], l3_line14[1], l3_line14[2], l2_line14[1], l2_line15[0]) ;

   FA level3_line15_FA1 ( l3_line15[0], l3_line15[1], l3_line15[2], l2_line15[1], l2_line16[0]) ;

   FA level3_line16_FA1 ( l3_line16[0], l3_line16[1], l3_line16[2], l2_line16[1], l2_line17[0]) ;

   FA level3_line17_FA1 ( l3_line17[0], l3_line17[1], l3_line17[2], l2_line17[1], l2_line18[0]) ;

   FA level3_line18_FA1 ( l3_line18[0], l3_line18[1], l3_line18[2], l2_line18[1], l2_line19[0]) ;

   FA level3_line19_FA1 ( l3_line19[0], l3_line19[1], l3_line19[2], l2_line19[1], l2_line20[0]) ;

   FA level3_line20_FA1 ( l3_line20[0], l3_line20[1], l3_line20[2], l2_line20[1], l2_line21[0]) ;

   FA level3_line21_FA1 ( l3_line21[0], l3_line21[1], l3_line21[2], l2_line21[1], l2_line22[0]) ;

   FA level3_line22_FA1 ( l3_line22[0], l3_line22[1], l3_line22[2], l2_line22[1], l2_line23[0]) ;

   FA level3_line23_FA1 ( l3_line23[0], l3_line23[1], l3_line23[2], l2_line23[1], l2_line24[0]) ;

   FA level3_line24_FA1 ( l3_line24[0], l3_line24[1], l3_line24[2], l2_line24[1], l2_line25[0]) ;

   FA level3_line25_FA1 ( l3_line25[0], l3_line25[1], l3_line25[2], l2_line25[1], l2_line26[0]) ;

   FA level3_line26_FA1 ( l3_line26[0], l3_line26[1], l3_line26[2], l2_line26[1], l2_line27[0]) ;

   FA level3_line27_FA1 ( l3_line27[0], l3_line27[1], l3_line27[2], l2_line27[1], l2_line28[0]) ;

   FA level3_line28_FA1 ( l3_line28[0], l3_line28[1], l3_line28[2], l2_line28[1], l2_line29[0]) ;

   FA level3_line29_FA1 ( l3_line29[0], l3_line29[1], l3_line29[2], l2_line29[1], l2_line30[0]) ;

   FA level3_line30_FA1 ( l3_line30[0], l3_line30[1], l3_line30[2], l2_line30[1], l2_line31[0]) ;

   FA level3_line31_FA1 ( l3_line31[0], l3_line31[1], l3_line31[2], l2_line31[1], l2_line32[0]) ;

   FA level3_line32_FA1 ( l3_line32[0], l3_line32[1], l3_line32[2], l2_line32[1], l2_line33[0]) ;

   FA level3_line33_FA1 ( l3_line33[0], l3_line33[1], l3_line33[2], l2_line33[1], l2_line34[0]) ;

   FA level3_line34_FA1 ( l3_line34[0], l3_line34[1], l3_line34[2], l2_line34[1], l2_line35[0]) ;

   FA level3_line35_FA1 ( l3_line35[0], l3_line35[1], l3_line35[2], l2_line35[1], l2_line36[0]) ;
	
	assign l2_line5[2] = l3_line5[3] ;
   assign l2_line6[2] = l3_line6[3] ;
   assign l2_line7[2] = l3_line7[3] ;
   assign l2_line8[2] = l3_line8[3] ;
   assign l2_line9[2] = l3_line9[3] ;
   assign l2_line10[2] = l3_line10[3] ;
   assign l2_line11[2] = l3_line11[3] ;
   assign l2_line12[2] = l3_line12[3] ;
   assign l2_line13[2] = l3_line13[3] ;
   assign l2_line14[2] = l3_line14[3] ;
   assign l2_line15[2] = l3_line15[3] ;
   assign l2_line16[2] = l3_line16[3] ;
   assign l2_line17[2] = l3_line17[3] ;
   assign l2_line18[2] = l3_line18[3] ;
   assign l2_line19[2] = l3_line19[3] ;
   assign l2_line20[2] = l3_line20[3] ;
   assign l2_line21[2] = l3_line21[3] ;
   assign l2_line22[2] = l3_line22[3] ;
   assign l2_line23[2] = l3_line23[3] ;
   assign l2_line24[2] = l3_line24[3] ;
   assign l2_line25[2] = l3_line25[3] ;
   assign l2_line26[2] = l3_line26[3] ;
   assign l2_line27[2] = l3_line27[3] ;
   assign l2_line28[2] = l3_line28[3] ;
   assign l2_line29[2] = l3_line29[3] ;
   assign l2_line30[2] = l3_line30[3] ;
   assign l2_line31[2] = l3_line31[3] ;
   assign l2_line32[2] = l3_line32[3] ;
   assign l2_line33[2] = l3_line33[3] ;
   assign l2_line34[2] = l3_line34[3] ;
   assign l2_line35[2] = l3_line35[3] ;
	assign l2_line36[2:1] = l3_line36[1:0] ;
	
	// passing first 3 level-3 lines as it is to nect level with capacity of 3 wires
	assign l2_line1 = l3_line1 ;
   assign l2_line2 = l3_line2 ;
   assign l2_line3 = l3_line3 ;
	
	//passing rest of the values which will be passed to next level as it is
   assign l2_line37 = l3_line37 ;
	
	// Level-3 (4) to level-2 (3) complete
	// Declaring level-1 lines
	wire       l1_line1 ;
	wire [1:0] l1_line2 ;
   wire [1:0] l1_line3 ;
   wire [1:0] l1_line4 ;
   wire [1:0] l1_line5 ;
   wire [1:0] l1_line6 ;
   wire [1:0] l1_line7 ;
   wire [1:0] l1_line8 ;
   wire [1:0] l1_line9 ;
   wire [1:0] l1_line10 ;
   wire [1:0] l1_line11 ;
   wire [1:0] l1_line12 ;
   wire [1:0] l1_line13 ;
   wire [1:0] l1_line14 ;
   wire [1:0] l1_line15 ;
   wire [1:0] l1_line16 ;
   wire [1:0] l1_line17 ;
   wire [1:0] l1_line18 ;
   wire [1:0] l1_line19 ;
   wire [1:0] l1_line20 ;
   wire [1:0] l1_line21 ;
   wire [1:0] l1_line22 ;
   wire [1:0] l1_line23 ;
   wire [1:0] l1_line24 ;
   wire [1:0] l1_line25 ;
   wire [1:0] l1_line26 ;
   wire [1:0] l1_line27 ;
   wire [1:0] l1_line28 ;
   wire [1:0] l1_line29 ;
   wire [1:0] l1_line30 ;
   wire [1:0] l1_line31 ;
   wire [1:0] l1_line32 ;
   wire [1:0] l1_line33 ;
   wire [1:0] l1_line34 ;
   wire [1:0] l1_line35 ;
   wire [1:0] l1_line36 ;
   wire [1:0] l1_line37 ;
	
	// passing first set of wires as it is
	assign l1_line1 = l2_line1 ;
	assign l1_line2 = l2_line2 ;
	
	// Full adder instantiation
	HA level2_line3_HA1 ( l2_line3[0], l2_line3[1],              l1_line3[0], l1_line4[0]) ;
	assign l1_line3[1] = l2_line3[2] ;
	
   FA level2_line4_FA1 ( l2_line4[0], l2_line4[1], l2_line4[2], l1_line4[1], l1_line5[0]) ;

   FA level2_line5_FA1 ( l2_line5[0], l2_line5[1], l2_line5[2], l1_line5[1], l1_line6[0]) ;

   FA level2_line6_FA1 ( l2_line6[0], l2_line6[1], l2_line6[2], l1_line6[1], l1_line7[0]) ;

   FA level2_line7_FA1 ( l2_line7[0], l2_line7[1], l2_line7[2], l1_line7[1], l1_line8[0]) ;

   FA level2_line8_FA1 ( l2_line8[0], l2_line8[1], l2_line8[2], l1_line8[1], l1_line9[0]) ;

   FA level2_line9_FA1 ( l2_line9[0], l2_line9[1], l2_line9[2], l1_line9[1], l1_line10[0]) ;

   FA level2_line10_FA1 ( l2_line10[0], l2_line10[1], l2_line10[2], l1_line10[1], l1_line11[0]) ;

   FA level2_line11_FA1 ( l2_line11[0], l2_line11[1], l2_line11[2], l1_line11[1], l1_line12[0]) ;

   FA level2_line12_FA1 ( l2_line12[0], l2_line12[1], l2_line12[2], l1_line12[1], l1_line13[0]) ;

   FA level2_line13_FA1 ( l2_line13[0], l2_line13[1], l2_line13[2], l1_line13[1], l1_line14[0]) ;

   FA level2_line14_FA1 ( l2_line14[0], l2_line14[1], l2_line14[2], l1_line14[1], l1_line15[0]) ;

   FA level2_line15_FA1 ( l2_line15[0], l2_line15[1], l2_line15[2], l1_line15[1], l1_line16[0]) ;

   FA level2_line16_FA1 ( l2_line16[0], l2_line16[1], l2_line16[2], l1_line16[1], l1_line17[0]) ;

   FA level2_line17_FA1 ( l2_line17[0], l2_line17[1], l2_line17[2], l1_line17[1], l1_line18[0]) ;

   FA level2_line18_FA1 ( l2_line18[0], l2_line18[1], l2_line18[2], l1_line18[1], l1_line19[0]) ;

   FA level2_line19_FA1 ( l2_line19[0], l2_line19[1], l2_line19[2], l1_line19[1], l1_line20[0]) ;

   FA level2_line20_FA1 ( l2_line20[0], l2_line20[1], l2_line20[2], l1_line20[1], l1_line21[0]) ;

   FA level2_line21_FA1 ( l2_line21[0], l2_line21[1], l2_line21[2], l1_line21[1], l1_line22[0]) ;

   FA level2_line22_FA1 ( l2_line22[0], l2_line22[1], l2_line22[2], l1_line22[1], l1_line23[0]) ;

   FA level2_line23_FA1 ( l2_line23[0], l2_line23[1], l2_line23[2], l1_line23[1], l1_line24[0]) ;

   FA level2_line24_FA1 ( l2_line24[0], l2_line24[1], l2_line24[2], l1_line24[1], l1_line25[0]) ;

   FA level2_line25_FA1 ( l2_line25[0], l2_line25[1], l2_line25[2], l1_line25[1], l1_line26[0]) ;

   FA level2_line26_FA1 ( l2_line26[0], l2_line26[1], l2_line26[2], l1_line26[1], l1_line27[0]) ;

   FA level2_line27_FA1 ( l2_line27[0], l2_line27[1], l2_line27[2], l1_line27[1], l1_line28[0]) ;

   FA level2_line28_FA1 ( l2_line28[0], l2_line28[1], l2_line28[2], l1_line28[1], l1_line29[0]) ;

   FA level2_line29_FA1 ( l2_line29[0], l2_line29[1], l2_line29[2], l1_line29[1], l1_line30[0]) ;

   FA level2_line30_FA1 ( l2_line30[0], l2_line30[1], l2_line30[2], l1_line30[1], l1_line31[0]) ;

   FA level2_line31_FA1 ( l2_line31[0], l2_line31[1], l2_line31[2], l1_line31[1], l1_line32[0]) ;

   FA level2_line32_FA1 ( l2_line32[0], l2_line32[1], l2_line32[2], l1_line32[1], l1_line33[0]) ;

   FA level2_line33_FA1 ( l2_line33[0], l2_line33[1], l2_line33[2], l1_line33[1], l1_line34[0]) ;

   FA level2_line34_FA1 ( l2_line34[0], l2_line34[1], l2_line34[2], l1_line34[1], l1_line35[0]) ;

   FA level2_line35_FA1 ( l2_line35[0], l2_line35[1], l2_line35[2], l1_line35[1], l1_line36[0]) ;

   FA level2_line36_FA1 ( l2_line36[0], l2_line36[1], l2_line36[2], l1_line36[1], l1_line37[0]) ;
	
	assign l1_line37[1] = l2_line37 ;
	
	wire [39:0] adder1_a,adder1_b ;// adder2_a,adder2_b ;
	wire adder1_cin; // adder2_cin ;
	wire [39:0] adder1_sum; // adder2_sum ;
	wire adder1_cout, adder2_cout ;
	
	assign adder1_cin = 1'b0 ;
	
	assign adder1_a[0] = 1'b0 ;//l1_line1[1] ;
   assign adder1_b[0] = l1_line1 ;
   assign adder1_a[1] = l1_line2[1] ;
   assign adder1_b[1] = l1_line2[0] ;
   assign adder1_a[2] = l1_line3[1] ;
   assign adder1_b[2] = l1_line3[0] ;
   assign adder1_a[3] = l1_line4[1] ;
   assign adder1_b[3] = l1_line4[0] ;
   assign adder1_a[4] = l1_line5[1] ;
   assign adder1_b[4] = l1_line5[0] ;
   assign adder1_a[5] = l1_line6[1] ;
   assign adder1_b[5] = l1_line6[0] ;
   assign adder1_a[6] = l1_line7[1] ;
   assign adder1_b[6] = l1_line7[0] ;
   assign adder1_a[7] = l1_line8[1] ;
   assign adder1_b[7] = l1_line8[0] ;
   assign adder1_a[8] = l1_line9[1] ;
   assign adder1_b[8] = l1_line9[0] ;
   assign adder1_a[9] = l1_line10[1] ;
   assign adder1_b[9] = l1_line10[0] ;
   assign adder1_a[10] = l1_line11[1] ;
   assign adder1_b[10] = l1_line11[0] ;
   assign adder1_a[11] = l1_line12[1] ;
   assign adder1_b[11] = l1_line12[0] ;
   assign adder1_a[12] = l1_line13[1] ;
   assign adder1_b[12] = l1_line13[0] ;
   assign adder1_a[13] = l1_line14[1] ;
   assign adder1_b[13] = l1_line14[0] ;
   assign adder1_a[14] = l1_line15[1] ;
   assign adder1_b[14] = l1_line15[0] ;
   assign adder1_a[15] = l1_line16[1] ;
   assign adder1_b[15] = l1_line16[0] ;
   assign adder1_a[16] = l1_line17[1] ;
   assign adder1_b[16] = l1_line17[0] ;
   assign adder1_a[17] = l1_line18[1] ;
   assign adder1_b[17] = l1_line18[0] ;
   assign adder1_a[18] = l1_line19[1] ;
   assign adder1_b[18] = l1_line19[0] ;
   assign adder1_a[19] = l1_line20[1] ;
   assign adder1_b[19] = l1_line20[0] ;
   assign adder1_a[20] = l1_line21[1] ;
   assign adder1_b[20] = l1_line21[0] ;
   assign adder1_a[21] = l1_line22[1] ;
   assign adder1_b[21] = l1_line22[0] ;
   assign adder1_a[22] = l1_line23[1] ;
   assign adder1_b[22] = l1_line23[0] ;
   assign adder1_a[23] = l1_line24[1] ;
   assign adder1_b[23] = l1_line24[0] ;
   assign adder1_a[24] = l1_line25[1] ;
   assign adder1_b[24] = l1_line25[0] ;
   assign adder1_a[25] = l1_line26[1] ;
   assign adder1_b[25] = l1_line26[0] ;
   assign adder1_a[26] = l1_line27[1] ;
   assign adder1_b[26] = l1_line27[0] ;
   assign adder1_a[27] = l1_line28[1] ;
   assign adder1_b[27] = l1_line28[0] ;
   assign adder1_a[28] = l1_line29[1] ;
   assign adder1_b[28] = l1_line29[0] ;
   assign adder1_a[29] = l1_line30[1] ;
   assign adder1_b[29] = l1_line30[0] ;
   assign adder1_a[30] = l1_line31[1] ;
   assign adder1_b[30] = l1_line31[0] ;
   assign adder1_a[31] = l1_line32[1] ;
   assign adder1_b[31] = l1_line32[0] ;
   assign adder1_a[32] = l1_line33[1] ;
   assign adder1_b[32] = l1_line33[0] ;
   assign adder1_a[33] = l1_line34[1] ;
   assign adder1_b[33] = l1_line34[0] ;
   assign adder1_a[34] = l1_line35[1] ;
   assign adder1_b[34] = l1_line35[0] ;
   assign adder1_a[35] = l1_line36[1] ;
   assign adder1_b[35] = l1_line36[0] ;
   assign adder1_a[36] = l1_line37[1] ;
   assign adder1_b[36] = l1_line37[0] ;
   assign adder1_a[37] = 1'b0 ;
   assign adder1_b[37] = 1'b0 ;
   assign adder1_a[38] = 1'b0 ;
   assign adder1_b[38] = 1'b0 ;
   assign adder1_a[39] = 1'b0 ;
   assign adder1_b[39] = 1'b0 ;
	
	adder_40_bit #(40) adder1 (adder1_a,adder1_b,adder1_cin,adder1_sum,adder1_cout) ;
	
	assign mul = adder1_sum[37:0] ;

endmodule
	